class apb_passive_agent_a2 extends uvm_agent;
  `uvm_component_utils(apb_passive_agent_a2)
  function new(string name="apb_passive_agent_a2",uvm_component parent);
    super.new(name,parent);
  endfunction
endclass
